`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 18.10.2022 22:02:00
// Design Name: 
// Module Name: FourDigitLEDdriver_testbench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module FourDigitLEDdriver_testbench;
    
    reg reset, clk;
    wire an3, an2, an1, an0;
    wire a, b, c, d, e, f, g, dp;
    
    
    
    
endmodule
